.param MOSFET_0_8_W_BIASCM_PMOS=5.2683098713337095 MOSFET_0_8_L_BIASCM_PMOS=0.8648659529510403 MOSFET_0_8_M_BIASCM_PMOS=42
.param MOSFET_8_2_W_gm1_PMOS=3.7458166970414863 MOSFET_8_2_L_gm1_PMOS=4.630555392006197 MOSFET_8_2_M_gm1_PMOS=13
.param MOSFET_10_1_W_gm2_PMOS=6.329021651180747 MOSFET_10_1_L_gm2_PMOS=3.9484141936873183 MOSFET_10_1_M_gm2_PMOS=46
.param MOSFET_11_1_W_gmf2_PMOS=4.693834488325472 MOSFET_11_1_L_gmf2_PMOS=0.7742450064609567 MOSFET_11_1_M_gmf2_PMOS=101
.param MOSFET_17_7_W_BIASCM_NMOS=1.00419582131841 MOSFET_17_7_L_BIASCM_NMOS=0.9347001989413464 MOSFET_17_7_M_BIASCM_NMOS=26
.param MOSFET_21_2_W_LOAD2_NMOS=5.871574021887089 MOSFET_21_2_L_LOAD2_NMOS=1.9200314285315998 MOSFET_21_2_M_LOAD2_NMOS=41
.param MOSFET_23_1_W_gm3_NMOS=0.792970207556583 MOSFET_23_1_L_gm3_NMOS=4.632315427792695 MOSFET_23_1_M_gm3_NMOS=30
.param CURRENT_0_BIAS=2.8539724202703217e-05
.param M_C0=19
.param M_C1=20
